module lifo #(
  parameter int DWIDTH        = 16,
  parameter int AWIDTH        = 8,
  parameter int ALMOST_FULL   = 2,
  parameter int ALMOST_EMPTY  = 2
)(
  input               clk_i,
  input               srst_i,

  input               wrreq_i,
  input  [DWIDTH-1:0] data_i,

  input               rdreq_i,
  output [DWIDTH-1:0] q_o,

  output              almost_empty_o,
  output              empty_o,
  output              almost_full_o,
  output              full_o,
  output [AWIDTH:0]   usedw_o
);

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "ModelSim" , encrypt_agent_info = "10.5b"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
kdexpbBKBPBuadRs2OKe4UdTznt7CSnNg4SGCh7B1uwBdWihKu6F9ntESfDRNnm2
A+Tv4Co/XUjW0jiXi6RH8cCIdDpPU/WKLYTvGo1R1ck6M/7jcNHRA+I4vnFIumim
OBPoUv4k+Fi0MIw2zP/rgZrGm8cF6WJXnNLyzpf4/NunyWVIu6td0g2T9ArhHUl2
pSJLBPx2SUgFivWOBKwIVt2bv8H6gYmT+Oz1YjiMVYMeN50+tDmjyGjn3noi725s
Pf1Oup5w+uNuwv4u0TZkztzM6iOb5dT4zkGVoJNfVyarq16fdNNWauKt2ZJwdfKs
spDqV79THVq1PAGLokF6cA==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 4528 )
`pragma protect data_block
FSXkNz6sODVCAb4YmmJ+sOkCMv3TU5PXAOC59ZHxsh3Xer8eeKlEYfOFlOL4mily
JijC25CtmvLJe2itWk+UVoN1Qjlvue3JrRjtWDEL5O5y6uUgbjWQlfjhSHqOJ+3f
J7TlK/nUYXpzUJsCgy0C5ODzA7D+js1wKVP/bdjwIEcTh/j5KEBG+FVjdoi6bRTe
r6GCdT57cGK8I1MjpEVs4xjrr47noQE5/cdYIYPz3PZHWAP0pf2gzp/RWpVhou2I
yJSVl09xP3rLHi02t6FhbiwXFSpA8SUS7V4ZDAW4zVA+Ome6kVoetEkQpUOc6fVf
zzoqCIWQ869lWVtT1lE599OvakAwE6zPuMacjD0Bt9M+Qeoypoq3PYkt455aKTuA
72HBLFxIDWs+uRzX8RMJpzMYCWpmlTPHwIXpFronLF5Tdesctd0mRjHY0Up3tUV/
hxfRpObCYUsqwFRKxWaG44qjS9kVvwHZlyu/zZKmvtXSJCuLhkAjEt0eOKew4LE7
9ResJgN6Z/QI71M03+08GvFuLtzu4SOvdkUFi7orgqqs4+HH34W7qpHlv5iQZNY0
Acl8yLQtYyjpM61+2g+cM0Lka4XoABswD1SlmTp8nxDlQLqkjcJhlppOKjqibgLV
69Fi2fdUHMiKDqyfZCYK7ABbHv3Aiw2ABvnoYLdDTbuGYgeq/EgJDvqToyz0R1CD
aRXkd05jLVbOBUQSRMiRSJKsI1cJRQe33v8QZZtwL6WrbfZVPfYYw7mKNzM30GbN
2IB5XrINOL4HBjfajF7Sp+075pRKU12MJnK2olWK7fTcVfH4qXsHtf2x6OjGaukR
dJBxbnUPiWPuUezK21R5BsMaCXy0anKWgx33kGvF24q3KinSFSWb9fMJbba2YPYe
x0PwyagZJu7JhPAwJ451JhYbV3H2xtkxJGX3Ac9rYp5H7X8YWP55wiaJ1yx53H0d
HOVwvGoOnMFg2yY4oWIO4vgLWfPnE1ZGwCREpU92jt8UmnmXKjYGXMIGeTdDKKbQ
MLbTReZlHpxxJR2Hxs2gz+ZXmQ3FZZzvZk2pyP5mTdcmDMEP32nuh/Tl8BTkDvld
V8My/UPxogLlCL+jMzjLqJh9hXpSZiTYtD+4JlD5zKHgLIRuNlq7an/zmt7F28mR
dHUPIj/TwkR0jfBEqYfmF/msFVC++kfA+xDcZYSICZAOgdHKYV91cZhnT35TBboH
i3hjMhIiAqqxm+J320t7lk5FpvJyN7iExVxW5DJl6v+NJqf0XlVXauX4Ca84FGGw
MorYlXxYExRnsvbkvleWSkB0GRfFAZfuTXwnSUew0H/hl7TgeYZxxcuthHUDKc6Q
huQxkmxs067YQ2C7D6pQ98GnkYSP8qUvRxAKZSMgHNSQP/GPOv39KDl1WhWq48p9
eRbMEnHHEhZBuQSzeVo/eDdyASeBizg1I034zdGJfVAvu4vUs9WD8qiJz6n5NrDY
l5QjK40Gm9ctVej3UvjZAJ9coX+gsINE7Z60kw+ZvVV/va4s537xR1X5kykeP4GH
zdUvKGK7X0q/C6Zcaa9ApoC3NCvF0f4A8Z6KOyzSDlrpQe5NDHaGwDHic8rlBSgR
FHqC6dpp0DmOrfcx7IL32O92V8f9iLk2ThlUAGSgzj9AYWCugMULsfN8KPMgDHWl
e+Py8kFhWrOg9UymFCTVYNLV9skemEhnojXd3tbriY/G9NpuhLwk+jbBxPuX9vBs
v+ALIkYEzePjotgwnr1OmNV2BHdWtAUT6E2KRvz9Qu5lWP5AKUk5VPIFDqDgVGIB
PIyNyM+Z2F4oZif9OZp/O9dWc350W+IZZOgACU4DoMqJfo6DHUWj2YWn5t1Ql7gy
TbsfaiHpqgqnVOiAJ0py820WDhERQE4SF5SaYd3XpMtLCtNOkXta+Bc8f/f7GIqQ
G/Or9fsG2IphfW1//9H2FpaeyTEwLFQJS5pzNHLPCSi4AHGUoxkEdD+FVCoylky5
vlziYUz67pgdEBIL/9pTXXV/Cf3scMf1uD+ClVw1vlCG58mSDeh4pLufojgW1o7a
s1cwWob2vmKzz1xzL34iDWxiwW2XMwd4gyLpXJkLSJTVlJo4BCK1lfOM/X8kHsz5
CTJsoYAZmOFi7ufXVI2v1uCznyRhAKokXhf2ZpNszw6MAN2aDWFLMHYrSz2xaTkX
MzfAYb22gFDJmo3ogi/QBOeJQbYgQdvASEBMNBhBHdz4ZGWktmDDuiu0p1Cki6wx
B4iBd4B/MQKPmanyub+EkwvFLO6ALGJqsrjCJlVskl0VTLHtFwmMy1OTxMDaa7O7
2c+HZWNsQREV+w79YxZrJBADrJkk2rHCGjQxdZE0YNLii3zvknOKR8p0nEOaiH/4
iXVCtluIhk7gA/LUwedJWfg+SB67a+NPZcFALCGFPary+YJYfQDg9XTKqi3K6AQd
GWxsoIMBFQRxGu/4JBilILf0Z6NgD5ZZAEU4TUVu0qcWcaK3btwuhjst0JbJbyD1
56Nro27W9q9Dxb5e73Vp/r6Xouq+8aSzQFYNVa8yDDJiYKMt7anfUBamARKmYJcL
osfdevlh0liBGaVUkmv9NxkdS4Bc1o04DaaJaUsmhCwC+T+PErD1T4GZq00cTgbi
XqLAMbkfc8Y+tqOwo3f2b0b3m60Ob6f8bY7Xsj54QE1RCjRsVbZszloAsxHEXPdx
e5oXx9a7FCqBVwWT0C68lakhAseSFqjvuKzNX3GfaA8bWJpNq4ciyE1km95D20sT
1imjcho09t4FiNzucSVv+BMzgo7wdiRBJi4iraXbiQBd/ORJ8OxSvsDXdcRlekNM
D7hshWFvBOovcHTphjIdlgfsFEVx1ozW7DagJ9YukZkmuzpS4cfso0z2HejdfZ3W
HiGM93ifk27w5gSwca8RZ1CMDdYulkj56/SqtLFBs2jBB/LrsEhwpQMWYLFvm0oG
MnaMV8zjtTiv66pR2H2owwS9Rnh6f4Pl4hsRDhOYbXx1GwJEFM6yZPQiNhJ/qWH2
JWrjTbriYMEVZ+9GAMV/v6CzqSMG4gW6MkjBKW+RvVZm6yD+5SiJ5z2dZ1s7PlCZ
jYBmwRX9I0zAAP9AdQH/miiXP1fRpEaPW48NbfZiccjwU72u+XYw1MpgMGn9xgKO
YYbC+L2SpXxKxg7IFgHBBfcc9bkLaQavkCiKiYIxSELP8WOd9KdxUiC2qYEOsAcM
g7mx4Zwss23sg7/h2AlsuwJmVxfr3OhgJqYSXPfed2XgscTU2w+RFGNebuF3spyC
Ij9a3tHVcJ0MSpdBRTfkLo5gnRr0EWoCECNaXge3hPVriVhEs3Y7OshAr5iEgvVP
Jab8rg5LypBqIv9KQ6jRCKxHuFGBphfPejEEZH1wreD87g18PHEYFkHaIcB92c9f
MMQi3a1r0qeePMq9i6TpXnwy4nhhBL09IxB/bkACHgDvdCOfcMcu3MfD1mntblKE
jo+zFqxQ96wNH+hh5wP1+XgxFLf9/SpIMIYaGKWGtVjueyMm+8ETHKloJ4yTiF/2
p3yJSiLaoW90eCS3F9Cm3kXG2hO9N80TTRSdbnCNUcy2xD1CpsGJf88EBjbKwKdV
TV05Fj3aOx/noCHzcdzRMXfzQGJa2QPqL+Wu27aGF9anQ3uap9PhbcAUvMVywLqk
WHUUQyDqr5HXU0RGpw3N2fLxBH1p8nLn0v6P7HrvPj5aRK/JK2ZVmDOEQ9k+ZjUa
GNW27T3oSqotuL9528Pf5hBK2eBf11BZmRMoG4CtWlKIeYXR/RjCZ441PiUuUWZs
x0nFd4eHqrveN/tm4RiFkGg8krdX5ozlQ1MQrYUn/V55RU4+u4zaGikvZsqhoRKk
LgsmRGFxTQPB2plnDf05qeiylrEayugb9PQPREu473t4eN6RBB6iUjwAteNKSejN
9MlNQEIyMf2sciVngrz+Ewy4fjQE4ZHXKlXaMUzf2r+6R7r0L0PugcUv3dvlw/07
ALEOH14poK4vhk7NSk4HBY3oX+NnviRittNolC6zp7hkFdGC0MdYWP3xy/LsmsU8
1pFitgL+WvDncT2wyB8HXFjwL0/bRL054DcmlLXHgGcVddkX0f/l3YNNX4AYi51G
tKNbKOlMW3H7FD3mOSUM0/HcUXrO/LqBwYw95uZBeo0jy/ktH5ExJfq6rZJMogLt
Y3MIysRulJFx3ClYId1lPmclVorjeO2id/DzTyUVa6/D2HizLU2TP2vEjiLhLFqY
67K+5CSpBOop8i4+jflc4sUq++JkXyepSuwdolntJVHwMB5pbosbM4lJCLfdun0w
B5Lx2cbxzydqRzppwRWRahm4oKOIEovUI/qcWktiGfu+42As8cWVa1VqleNaEpmp
dsxhbYB+IyskWJPo9LSH3MTWe6K1ELuiNtTnxALZF/+XOTSFZck21PoeOpXYuEQf
ayvaeOCgGyK+g/D1r9C/Hh4ewkiBj3L5gLBpnEGmCFW3+yMNUNqWH0WzU5E0vEwV
hgF5zJ63vLiVciOqZPl2hywXnTzHbJrA6BtLpeH9gLmlVQ5zTxsGwzUzFsYoYSlK
a6fp26elEmAPlmufO3iUY8TVirAf30Wkm5i9ir74+zV3rfMoN7S0CCZ0goqM3Muw
vht1pkbvrf68dlFQKscSqy4PXe9YBbodBVAnwEeWxh78SOPAYNu+fU0QZ52RdtmU
B06nV8d84jDbdpb8tDPbr31VShqYP4YYFodhA12D5kXh8rWb2vARdz6xq5E+neEr
P3TY4sJQFZdSOcGiUaT8rHHyiRC0NGylM17SQJyrkLA1vSgfhyPG18dIbVd3SuYo
aacpr0EffI6uBTv6XTrs/VLCNSq8qp86kckwaURZL+8uPpqLB11n2S4uIdJH63Xb
U++sp37fvzW3aov3eQ2o4onjluos6+i0ovy0JCXfiMBYPUCHhiY2oABPrRdWQn5G
tHDiMFaRfgBBS62kYPAUXdJ2RF+DqCIJ5aBJOJgdnXmcG2vn6qWKeQEH+vHbmcJz
kWCdjkkqpV8tUQCF99ny3CdlYN+KmAQ/3hPN+eYb3WnhZCt+jhvrIaZW/e0kKfok
7cZqrvadV9r9NKlJ6d2jEexlkyM4DB9lLuvqr7db/x7L4JObCYFnUH+zdqIGVC2S
ho9+o+x2wnWJGBTRjng2wbTaCTBcR//27hcBRtEwCrvUitbL+8fRfue33BI/JfVj
46Xt1Wf+3fRdy79NnFloFaoaTkJG4uztMWZjg1mUr8uvTEPGbCB40bPfj7fWo5L5
DzKABiIQmdZlCuaTMMCgEio+4O1ZqOnBZOAD5EYMKur6fl3X4178F9Warm1Y2A5u
DCOTYJzTlzYs5DqTEQfURxO4v++hCSocwl+egp9YV17O1Z4zYGmdMHAufNzmXMD1
6zmT4b0+pdBPBS+9B6nmnjE3Uy0GZyG9kJlYHiR5KdBBpbvRrydtvJ1APBsDwRxr
ZW/KXrbEjFy9ZsxLNgdXw0DLHkXSFNf2S5P3euNt5m0X35n0fcGmeS+NDGsEvy6i
q7f3wvJK+klM5HalR+npdzpXjy9IBpZDXcL1lHTaSg0oLM594gA0QbLuq6gALrpr
p/CJf5slq9aHDYn2n+SHLKCfnrUGr46Trpsh0Dc6vNVLu9sezuOjgh6FjIycQWn7
ltcXqwI/ZkfB+SgwVH+K8RUXkR4As9/hqpuMOdEUFh4kjlVK1yRzN2PZWyiQRsB6
XI39wOiFgI1I4B0MqP2IFdjpJ2aTiB1eWUm+0WqnoeXKWQXrhU9LD992TpDXbWJB
jPetOk486SJMk0mfGEBmInol+NnzdMvdSUsqfXvurly2qYPmHXdmieyvhUtYXwMW
UL7bGV2ofLMpLBXbNY6sroL2ui0fQ5u5ErFUiFxIGhCZxj/6Kz9tFwtBbkITzxnn
Xcm0q2+tlZn57Jo5YJrS0RZo+FokPLH+eNve5NveqQPfu9Z2Dmhiv95bn5Kk7H8w
9NEdZF8WdCP22ethcdR0B/eJO4C2J7b3/TW4vjkVxbOAOA7C1KBFdvRXGIOCUKAL
Z82Kg2BOWHluA3FPMr5QLw==
`pragma protect end_protected
