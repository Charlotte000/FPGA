package byte_inc_package;

`include "byte_inc/byte_inc_transaction.sv"

`include "byte_inc/byte_inc_driver.sv"
`include "byte_inc/byte_inc_monitor.sv"
`include "byte_inc/byte_inc_agent.sv"

`include "byte_inc_generator.sv"
`include "byte_inc_scoreboard.sv"
`include "byte_inc_environment.sv"

endpackage
