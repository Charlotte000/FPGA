module bit_population_counter #(
  parameter int unsigned WIDTH,
  parameter int unsigned PIPELINE_SIZE
)(
  input  logic                   clk_i,
  input  logic                   srst_i,

  input  logic [WIDTH-1:0]       data_i,
  input  logic                   data_val_i,

  output logic [$clog2(WIDTH):0] data_o,
  output logic                   data_val_o
);

localparam int unsigned PIPELINE_COUNT = ( WIDTH / PIPELINE_SIZE );

logic [PIPELINE_COUNT:0][WIDTH-1:0]       pipeline_data;
logic [PIPELINE_COUNT:0]                  pipeline_data_val;
logic [PIPELINE_COUNT:0][$clog2(WIDTH):0] pipeline_count;

genvar i;
generate
  for( i = 0; i < PIPELINE_COUNT; i++ )
    begin : pipeline_generator
      bit_counter_pipeline #(
        .WIDTH           ( WIDTH             ),
        .PIPELINE_SIZE   ( PIPELINE_SIZE     ),
        .PIPELINE_OFFSET ( i * PIPELINE_SIZE )
      ) bit_counter_pipeline_inst (
        .clk_i      ( clk_i                  ),
        .data_i     ( pipeline_data[i]       ),
        .data_val_i ( pipeline_data_val[i]   ),
        .count_i    ( pipeline_count[i]      ),
        .data_o     ( pipeline_data[i+1]     ),
        .data_val_o ( pipeline_data_val[i+1] ),
        .count_o    ( pipeline_count[i+1]    )
      );
    end
endgenerate

always_ff @( posedge clk_i )
  pipeline_data[0] <= data_i;

always_ff @( posedge clk_i )
  pipeline_data_val[0] <= data_val_i;

always_ff @( posedge clk_i )
  data_o <= pipeline_count[PIPELINE_COUNT];

always_ff @( posedge clk_i )
  data_val_o <= pipeline_data_val[PIPELINE_COUNT];

assign pipeline_count[0] = '0;

endmodule
