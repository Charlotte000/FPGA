package ast_dmx_package;

`include "ast_dmx_packet.sv"

`include "ast_dmx_generator.sv"
`include "ast_dmx_driver.sv"
`include "ast_dmx_monitor.sv"
`include "ast_dmx_scoreboard.sv"
`include "ast_dmx_environment.sv"

endpackage
